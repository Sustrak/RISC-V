-- AvalonMM.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity AvalonMM is
	port (
		clk_clk                   : in    std_logic                     := '0';             --         clk.clk
		mm_bridge_s_waitrequest   : out   std_logic;                                        -- mm_bridge_s.waitrequest
		mm_bridge_s_readdata      : out   std_logic_vector(31 downto 0);                    --            .readdata
		mm_bridge_s_readdatavalid : out   std_logic;                                        --            .readdatavalid
		mm_bridge_s_burstcount    : in    std_logic_vector(0 downto 0)  := (others => '0'); --            .burstcount
		mm_bridge_s_writedata     : in    std_logic_vector(31 downto 0) := (others => '0'); --            .writedata
		mm_bridge_s_address       : in    std_logic_vector(27 downto 0) := (others => '0'); --            .address
		mm_bridge_s_write         : in    std_logic                     := '0';             --            .write
		mm_bridge_s_read          : in    std_logic                     := '0';             --            .read
		mm_bridge_s_byteenable    : in    std_logic_vector(3 downto 0)  := (others => '0'); --            .byteenable
		mm_bridge_s_debugaccess   : in    std_logic                     := '0';             --            .debugaccess
		pp_hex_03_HEX0            : out   std_logic_vector(6 downto 0);                     --   pp_hex_03.HEX0
		pp_hex_03_HEX1            : out   std_logic_vector(6 downto 0);                     --            .HEX1
		pp_hex_03_HEX2            : out   std_logic_vector(6 downto 0);                     --            .HEX2
		pp_hex_03_HEX3            : out   std_logic_vector(6 downto 0);                     --            .HEX3
		pp_hex_47_HEX4            : out   std_logic_vector(6 downto 0);                     --   pp_hex_47.HEX4
		pp_hex_47_HEX5            : out   std_logic_vector(6 downto 0);                     --            .HEX5
		pp_hex_47_HEX6            : out   std_logic_vector(6 downto 0);                     --            .HEX6
		pp_hex_47_HEX7            : out   std_logic_vector(6 downto 0);                     --            .HEX7
		pp_key_export             : in    std_logic_vector(3 downto 0)  := (others => '0'); --      pp_key.export
		pp_led_g_export           : out   std_logic_vector(8 downto 0);                     --    pp_led_g.export
		pp_led_r_export           : out   std_logic_vector(17 downto 0);                    --    pp_led_r.export
		pp_switch_export          : in    std_logic_vector(17 downto 0) := (others => '0'); --   pp_switch.export
		reset_reset_n             : in    std_logic                     := '0';             --       reset.reset_n
		sdram_addr                : out   std_logic_vector(12 downto 0);                    --       sdram.addr
		sdram_ba                  : out   std_logic_vector(1 downto 0);                     --            .ba
		sdram_cas_n               : out   std_logic;                                        --            .cas_n
		sdram_cke                 : out   std_logic;                                        --            .cke
		sdram_cs_n                : out   std_logic;                                        --            .cs_n
		sdram_dq                  : inout std_logic_vector(31 downto 0) := (others => '0'); --            .dq
		sdram_dqm                 : out   std_logic_vector(3 downto 0);                     --            .dqm
		sdram_ras_n               : out   std_logic;                                        --            .ras_n
		sdram_we_n                : out   std_logic;                                        --            .we_n
		sdram_clk_clk             : out   std_logic;                                        --   sdram_clk.clk
		switch_int_irq            : out   std_logic                                         --  switch_int.irq
	);
end entity AvalonMM;

architecture rtl of AvalonMM is
	component AvalonMM_hex_03 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			HEX0       : out std_logic_vector(6 downto 0);                     -- export
			HEX1       : out std_logic_vector(6 downto 0);                     -- export
			HEX2       : out std_logic_vector(6 downto 0);                     -- export
			HEX3       : out std_logic_vector(6 downto 0)                      -- export
		);
	end component AvalonMM_hex_03;

	component AvalonMM_hex_47 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			HEX4       : out std_logic_vector(6 downto 0);                     -- export
			HEX5       : out std_logic_vector(6 downto 0);                     -- export
			HEX6       : out std_logic_vector(6 downto 0);                     -- export
			HEX7       : out std_logic_vector(6 downto 0)                      -- export
		);
	end component AvalonMM_hex_47;

	component AvalonMM_jtag_master is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component AvalonMM_jtag_master;

	component AvalonMM_key is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			KEY        : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component AvalonMM_key;

	component AvalonMM_led_g is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			LEDG       : out std_logic_vector(8 downto 0)                      -- export
		);
	end component AvalonMM_led_g;

	component AvalonMM_led_r is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			LEDR       : out std_logic_vector(17 downto 0)                     -- export
		);
	end component AvalonMM_led_r;

	component altera_avalon_mm_bridge is
		generic (
			DATA_WIDTH        : integer := 32;
			SYMBOL_WIDTH      : integer := 8;
			HDL_ADDR_WIDTH    : integer := 10;
			BURSTCOUNT_WIDTH  : integer := 1;
			PIPELINE_COMMAND  : integer := 1;
			PIPELINE_RESPONSE : integer := 1
		);
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(27 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic;                                        -- debugaccess
			s0_response      : out std_logic_vector(1 downto 0);                     -- response
			m0_response      : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- response
		);
	end component altera_avalon_mm_bridge;

	component AvalonMM_sdram_controller is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(31 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(31 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(3 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component AvalonMM_sdram_controller;

	component AvalonMM_sdram_pll is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component AvalonMM_sdram_pll;

	component AvalonMM_switch is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			SW         : in  std_logic_vector(17 downto 0) := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component AvalonMM_switch;

	component AvalonMM_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                      : in  std_logic                     := 'X';             -- clk
			sdram_pll_sys_clk_clk                              : in  std_logic                     := 'X';             -- clk
			jtag_master_clk_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			led_r_reset_reset_bridge_in_reset_reset            : in  std_logic                     := 'X';             -- reset
			mm_bridge_reset_reset_bridge_in_reset_reset        : in  std_logic                     := 'X';             -- reset
			sdram_controller_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			jtag_master_master_address                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			jtag_master_master_waitrequest                     : out std_logic;                                        -- waitrequest
			jtag_master_master_byteenable                      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_master_master_read                            : in  std_logic                     := 'X';             -- read
			jtag_master_master_readdata                        : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_master_master_readdatavalid                   : out std_logic;                                        -- readdatavalid
			jtag_master_master_write                           : in  std_logic                     := 'X';             -- write
			jtag_master_master_writedata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			mm_bridge_m0_address                               : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			mm_bridge_m0_waitrequest                           : out std_logic;                                        -- waitrequest
			mm_bridge_m0_burstcount                            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			mm_bridge_m0_byteenable                            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			mm_bridge_m0_read                                  : in  std_logic                     := 'X';             -- read
			mm_bridge_m0_readdata                              : out std_logic_vector(31 downto 0);                    -- readdata
			mm_bridge_m0_readdatavalid                         : out std_logic;                                        -- readdatavalid
			mm_bridge_m0_write                                 : in  std_logic                     := 'X';             -- write
			mm_bridge_m0_writedata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			mm_bridge_m0_debugaccess                           : in  std_logic                     := 'X';             -- debugaccess
			hex_03_avalon_parallel_port_slave_address          : out std_logic_vector(1 downto 0);                     -- address
			hex_03_avalon_parallel_port_slave_write            : out std_logic;                                        -- write
			hex_03_avalon_parallel_port_slave_read             : out std_logic;                                        -- read
			hex_03_avalon_parallel_port_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex_03_avalon_parallel_port_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			hex_03_avalon_parallel_port_slave_byteenable       : out std_logic_vector(3 downto 0);                     -- byteenable
			hex_03_avalon_parallel_port_slave_chipselect       : out std_logic;                                        -- chipselect
			hex_47_avalon_parallel_port_slave_address          : out std_logic_vector(1 downto 0);                     -- address
			hex_47_avalon_parallel_port_slave_write            : out std_logic;                                        -- write
			hex_47_avalon_parallel_port_slave_read             : out std_logic;                                        -- read
			hex_47_avalon_parallel_port_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex_47_avalon_parallel_port_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			hex_47_avalon_parallel_port_slave_byteenable       : out std_logic_vector(3 downto 0);                     -- byteenable
			hex_47_avalon_parallel_port_slave_chipselect       : out std_logic;                                        -- chipselect
			key_avalon_parallel_port_slave_address             : out std_logic_vector(1 downto 0);                     -- address
			key_avalon_parallel_port_slave_write               : out std_logic;                                        -- write
			key_avalon_parallel_port_slave_read                : out std_logic;                                        -- read
			key_avalon_parallel_port_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			key_avalon_parallel_port_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			key_avalon_parallel_port_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			key_avalon_parallel_port_slave_chipselect          : out std_logic;                                        -- chipselect
			led_g_avalon_parallel_port_slave_address           : out std_logic_vector(1 downto 0);                     -- address
			led_g_avalon_parallel_port_slave_write             : out std_logic;                                        -- write
			led_g_avalon_parallel_port_slave_read              : out std_logic;                                        -- read
			led_g_avalon_parallel_port_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_g_avalon_parallel_port_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			led_g_avalon_parallel_port_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			led_g_avalon_parallel_port_slave_chipselect        : out std_logic;                                        -- chipselect
			led_r_avalon_parallel_port_slave_address           : out std_logic_vector(1 downto 0);                     -- address
			led_r_avalon_parallel_port_slave_write             : out std_logic;                                        -- write
			led_r_avalon_parallel_port_slave_read              : out std_logic;                                        -- read
			led_r_avalon_parallel_port_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_r_avalon_parallel_port_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			led_r_avalon_parallel_port_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			led_r_avalon_parallel_port_slave_chipselect        : out std_logic;                                        -- chipselect
			sdram_controller_s1_address                        : out std_logic_vector(24 downto 0);                    -- address
			sdram_controller_s1_write                          : out std_logic;                                        -- write
			sdram_controller_s1_read                           : out std_logic;                                        -- read
			sdram_controller_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sdram_controller_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			sdram_controller_s1_byteenable                     : out std_logic_vector(3 downto 0);                     -- byteenable
			sdram_controller_s1_readdatavalid                  : in  std_logic                     := 'X';             -- readdatavalid
			sdram_controller_s1_waitrequest                    : in  std_logic                     := 'X';             -- waitrequest
			sdram_controller_s1_chipselect                     : out std_logic;                                        -- chipselect
			switch_avalon_parallel_port_slave_address          : out std_logic_vector(1 downto 0);                     -- address
			switch_avalon_parallel_port_slave_write            : out std_logic;                                        -- write
			switch_avalon_parallel_port_slave_read             : out std_logic;                                        -- read
			switch_avalon_parallel_port_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			switch_avalon_parallel_port_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			switch_avalon_parallel_port_slave_byteenable       : out std_logic_vector(3 downto 0);                     -- byteenable
			switch_avalon_parallel_port_slave_chipselect       : out std_logic                                         -- chipselect
		);
	end component AvalonMM_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal sdram_pll_sys_clk_clk                                          : std_logic;                     -- sdram_pll:sys_clk_clk -> [jtag_master:clk_clk, mm_bridge:clk, mm_interconnect_0:sdram_pll_sys_clk_clk, rst_controller_001:clk, rst_controller_002:clk, sdram_controller:clk]
	signal sdram_pll_reset_source_reset                                   : std_logic;                     -- sdram_pll:reset_source_reset -> [jtag_master:clk_reset_reset, rst_controller_001:reset_in0]
	signal mm_bridge_m0_waitrequest                                       : std_logic;                     -- mm_interconnect_0:mm_bridge_m0_waitrequest -> mm_bridge:m0_waitrequest
	signal mm_bridge_m0_readdata                                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:mm_bridge_m0_readdata -> mm_bridge:m0_readdata
	signal mm_bridge_m0_debugaccess                                       : std_logic;                     -- mm_bridge:m0_debugaccess -> mm_interconnect_0:mm_bridge_m0_debugaccess
	signal mm_bridge_m0_address                                           : std_logic_vector(27 downto 0); -- mm_bridge:m0_address -> mm_interconnect_0:mm_bridge_m0_address
	signal mm_bridge_m0_read                                              : std_logic;                     -- mm_bridge:m0_read -> mm_interconnect_0:mm_bridge_m0_read
	signal mm_bridge_m0_byteenable                                        : std_logic_vector(3 downto 0);  -- mm_bridge:m0_byteenable -> mm_interconnect_0:mm_bridge_m0_byteenable
	signal mm_bridge_m0_readdatavalid                                     : std_logic;                     -- mm_interconnect_0:mm_bridge_m0_readdatavalid -> mm_bridge:m0_readdatavalid
	signal mm_bridge_m0_writedata                                         : std_logic_vector(31 downto 0); -- mm_bridge:m0_writedata -> mm_interconnect_0:mm_bridge_m0_writedata
	signal mm_bridge_m0_write                                             : std_logic;                     -- mm_bridge:m0_write -> mm_interconnect_0:mm_bridge_m0_write
	signal mm_bridge_m0_burstcount                                        : std_logic_vector(0 downto 0);  -- mm_bridge:m0_burstcount -> mm_interconnect_0:mm_bridge_m0_burstcount
	signal jtag_master_master_readdata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_master_master_readdata -> jtag_master:master_readdata
	signal jtag_master_master_waitrequest                                 : std_logic;                     -- mm_interconnect_0:jtag_master_master_waitrequest -> jtag_master:master_waitrequest
	signal jtag_master_master_address                                     : std_logic_vector(31 downto 0); -- jtag_master:master_address -> mm_interconnect_0:jtag_master_master_address
	signal jtag_master_master_read                                        : std_logic;                     -- jtag_master:master_read -> mm_interconnect_0:jtag_master_master_read
	signal jtag_master_master_byteenable                                  : std_logic_vector(3 downto 0);  -- jtag_master:master_byteenable -> mm_interconnect_0:jtag_master_master_byteenable
	signal jtag_master_master_readdatavalid                               : std_logic;                     -- mm_interconnect_0:jtag_master_master_readdatavalid -> jtag_master:master_readdatavalid
	signal jtag_master_master_write                                       : std_logic;                     -- jtag_master:master_write -> mm_interconnect_0:jtag_master_master_write
	signal jtag_master_master_writedata                                   : std_logic_vector(31 downto 0); -- jtag_master:master_writedata -> mm_interconnect_0:jtag_master_master_writedata
	signal mm_interconnect_0_led_r_avalon_parallel_port_slave_chipselect  : std_logic;                     -- mm_interconnect_0:led_r_avalon_parallel_port_slave_chipselect -> led_r:chipselect
	signal mm_interconnect_0_led_r_avalon_parallel_port_slave_readdata    : std_logic_vector(31 downto 0); -- led_r:readdata -> mm_interconnect_0:led_r_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_led_r_avalon_parallel_port_slave_address     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_r_avalon_parallel_port_slave_address -> led_r:address
	signal mm_interconnect_0_led_r_avalon_parallel_port_slave_read        : std_logic;                     -- mm_interconnect_0:led_r_avalon_parallel_port_slave_read -> led_r:read
	signal mm_interconnect_0_led_r_avalon_parallel_port_slave_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:led_r_avalon_parallel_port_slave_byteenable -> led_r:byteenable
	signal mm_interconnect_0_led_r_avalon_parallel_port_slave_write       : std_logic;                     -- mm_interconnect_0:led_r_avalon_parallel_port_slave_write -> led_r:write
	signal mm_interconnect_0_led_r_avalon_parallel_port_slave_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_r_avalon_parallel_port_slave_writedata -> led_r:writedata
	signal mm_interconnect_0_hex_03_avalon_parallel_port_slave_chipselect : std_logic;                     -- mm_interconnect_0:hex_03_avalon_parallel_port_slave_chipselect -> hex_03:chipselect
	signal mm_interconnect_0_hex_03_avalon_parallel_port_slave_readdata   : std_logic_vector(31 downto 0); -- hex_03:readdata -> mm_interconnect_0:hex_03_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_hex_03_avalon_parallel_port_slave_address    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex_03_avalon_parallel_port_slave_address -> hex_03:address
	signal mm_interconnect_0_hex_03_avalon_parallel_port_slave_read       : std_logic;                     -- mm_interconnect_0:hex_03_avalon_parallel_port_slave_read -> hex_03:read
	signal mm_interconnect_0_hex_03_avalon_parallel_port_slave_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_0:hex_03_avalon_parallel_port_slave_byteenable -> hex_03:byteenable
	signal mm_interconnect_0_hex_03_avalon_parallel_port_slave_write      : std_logic;                     -- mm_interconnect_0:hex_03_avalon_parallel_port_slave_write -> hex_03:write
	signal mm_interconnect_0_hex_03_avalon_parallel_port_slave_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex_03_avalon_parallel_port_slave_writedata -> hex_03:writedata
	signal mm_interconnect_0_hex_47_avalon_parallel_port_slave_chipselect : std_logic;                     -- mm_interconnect_0:hex_47_avalon_parallel_port_slave_chipselect -> hex_47:chipselect
	signal mm_interconnect_0_hex_47_avalon_parallel_port_slave_readdata   : std_logic_vector(31 downto 0); -- hex_47:readdata -> mm_interconnect_0:hex_47_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_hex_47_avalon_parallel_port_slave_address    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex_47_avalon_parallel_port_slave_address -> hex_47:address
	signal mm_interconnect_0_hex_47_avalon_parallel_port_slave_read       : std_logic;                     -- mm_interconnect_0:hex_47_avalon_parallel_port_slave_read -> hex_47:read
	signal mm_interconnect_0_hex_47_avalon_parallel_port_slave_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_0:hex_47_avalon_parallel_port_slave_byteenable -> hex_47:byteenable
	signal mm_interconnect_0_hex_47_avalon_parallel_port_slave_write      : std_logic;                     -- mm_interconnect_0:hex_47_avalon_parallel_port_slave_write -> hex_47:write
	signal mm_interconnect_0_hex_47_avalon_parallel_port_slave_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex_47_avalon_parallel_port_slave_writedata -> hex_47:writedata
	signal mm_interconnect_0_key_avalon_parallel_port_slave_chipselect    : std_logic;                     -- mm_interconnect_0:key_avalon_parallel_port_slave_chipselect -> key:chipselect
	signal mm_interconnect_0_key_avalon_parallel_port_slave_readdata      : std_logic_vector(31 downto 0); -- key:readdata -> mm_interconnect_0:key_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_key_avalon_parallel_port_slave_address       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:key_avalon_parallel_port_slave_address -> key:address
	signal mm_interconnect_0_key_avalon_parallel_port_slave_read          : std_logic;                     -- mm_interconnect_0:key_avalon_parallel_port_slave_read -> key:read
	signal mm_interconnect_0_key_avalon_parallel_port_slave_byteenable    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:key_avalon_parallel_port_slave_byteenable -> key:byteenable
	signal mm_interconnect_0_key_avalon_parallel_port_slave_write         : std_logic;                     -- mm_interconnect_0:key_avalon_parallel_port_slave_write -> key:write
	signal mm_interconnect_0_key_avalon_parallel_port_slave_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:key_avalon_parallel_port_slave_writedata -> key:writedata
	signal mm_interconnect_0_switch_avalon_parallel_port_slave_chipselect : std_logic;                     -- mm_interconnect_0:switch_avalon_parallel_port_slave_chipselect -> switch:chipselect
	signal mm_interconnect_0_switch_avalon_parallel_port_slave_readdata   : std_logic_vector(31 downto 0); -- switch:readdata -> mm_interconnect_0:switch_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_switch_avalon_parallel_port_slave_address    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switch_avalon_parallel_port_slave_address -> switch:address
	signal mm_interconnect_0_switch_avalon_parallel_port_slave_read       : std_logic;                     -- mm_interconnect_0:switch_avalon_parallel_port_slave_read -> switch:read
	signal mm_interconnect_0_switch_avalon_parallel_port_slave_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_0:switch_avalon_parallel_port_slave_byteenable -> switch:byteenable
	signal mm_interconnect_0_switch_avalon_parallel_port_slave_write      : std_logic;                     -- mm_interconnect_0:switch_avalon_parallel_port_slave_write -> switch:write
	signal mm_interconnect_0_switch_avalon_parallel_port_slave_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:switch_avalon_parallel_port_slave_writedata -> switch:writedata
	signal mm_interconnect_0_led_g_avalon_parallel_port_slave_chipselect  : std_logic;                     -- mm_interconnect_0:led_g_avalon_parallel_port_slave_chipselect -> led_g:chipselect
	signal mm_interconnect_0_led_g_avalon_parallel_port_slave_readdata    : std_logic_vector(31 downto 0); -- led_g:readdata -> mm_interconnect_0:led_g_avalon_parallel_port_slave_readdata
	signal mm_interconnect_0_led_g_avalon_parallel_port_slave_address     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_g_avalon_parallel_port_slave_address -> led_g:address
	signal mm_interconnect_0_led_g_avalon_parallel_port_slave_read        : std_logic;                     -- mm_interconnect_0:led_g_avalon_parallel_port_slave_read -> led_g:read
	signal mm_interconnect_0_led_g_avalon_parallel_port_slave_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:led_g_avalon_parallel_port_slave_byteenable -> led_g:byteenable
	signal mm_interconnect_0_led_g_avalon_parallel_port_slave_write       : std_logic;                     -- mm_interconnect_0:led_g_avalon_parallel_port_slave_write -> led_g:write
	signal mm_interconnect_0_led_g_avalon_parallel_port_slave_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_g_avalon_parallel_port_slave_writedata -> led_g:writedata
	signal mm_interconnect_0_sdram_controller_s1_chipselect               : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	signal mm_interconnect_0_sdram_controller_s1_readdata                 : std_logic_vector(31 downto 0); -- sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	signal mm_interconnect_0_sdram_controller_s1_waitrequest              : std_logic;                     -- sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	signal mm_interconnect_0_sdram_controller_s1_address                  : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	signal mm_interconnect_0_sdram_controller_s1_read                     : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_read -> mm_interconnect_0_sdram_controller_s1_read:in
	signal mm_interconnect_0_sdram_controller_s1_byteenable               : std_logic_vector(3 downto 0);  -- mm_interconnect_0:sdram_controller_s1_byteenable -> mm_interconnect_0_sdram_controller_s1_byteenable:in
	signal mm_interconnect_0_sdram_controller_s1_readdatavalid            : std_logic;                     -- sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	signal mm_interconnect_0_sdram_controller_s1_write                    : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_write -> mm_interconnect_0_sdram_controller_s1_write:in
	signal mm_interconnect_0_sdram_controller_s1_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	signal rst_controller_reset_out_reset                                 : std_logic;                     -- rst_controller:reset_out -> [hex_03:reset, hex_47:reset, key:reset, led_g:reset, led_r:reset, mm_interconnect_0:led_r_reset_reset_bridge_in_reset_reset, sdram_pll:ref_reset_reset, switch:reset]
	signal rst_controller_001_reset_out_reset                             : std_logic;                     -- rst_controller_001:reset_out -> [mm_bridge:reset, mm_interconnect_0:jtag_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:mm_bridge_reset_reset_bridge_in_reset_reset]
	signal rst_controller_002_reset_out_reset                             : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:sdram_controller_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in]
	signal jtag_master_master_reset_reset                                 : std_logic;                     -- jtag_master:master_reset_reset -> rst_controller_002:reset_in0
	signal reset_reset_n_ports_inv                                        : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_sdram_controller_s1_read_ports_inv           : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_read:inv -> sdram_controller:az_rd_n
	signal mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv     : std_logic_vector(3 downto 0);  -- mm_interconnect_0_sdram_controller_s1_byteenable:inv -> sdram_controller:az_be_n
	signal mm_interconnect_0_sdram_controller_s1_write_ports_inv          : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_write:inv -> sdram_controller:az_wr_n
	signal rst_controller_002_reset_out_reset_ports_inv                   : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> sdram_controller:reset_n

begin

	hex_03 : component AvalonMM_hex_03
		port map (
			clk        => clk_clk,                                                        --                        clk.clk
			reset      => rst_controller_reset_out_reset,                                 --                      reset.reset
			address    => mm_interconnect_0_hex_03_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_hex_03_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_hex_03_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_hex_03_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_hex_03_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_hex_03_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_hex_03_avalon_parallel_port_slave_readdata,   --                           .readdata
			HEX0       => pp_hex_03_HEX0,                                                 --         external_interface.export
			HEX1       => pp_hex_03_HEX1,                                                 --                           .export
			HEX2       => pp_hex_03_HEX2,                                                 --                           .export
			HEX3       => pp_hex_03_HEX3                                                  --                           .export
		);

	hex_47 : component AvalonMM_hex_47
		port map (
			clk        => clk_clk,                                                        --                        clk.clk
			reset      => rst_controller_reset_out_reset,                                 --                      reset.reset
			address    => mm_interconnect_0_hex_47_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_hex_47_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_hex_47_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_hex_47_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_hex_47_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_hex_47_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_hex_47_avalon_parallel_port_slave_readdata,   --                           .readdata
			HEX4       => pp_hex_47_HEX4,                                                 --         external_interface.export
			HEX5       => pp_hex_47_HEX5,                                                 --                           .export
			HEX6       => pp_hex_47_HEX6,                                                 --                           .export
			HEX7       => pp_hex_47_HEX7                                                  --                           .export
		);

	jtag_master : component AvalonMM_jtag_master
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => sdram_pll_sys_clk_clk,            --          clk.clk
			clk_reset_reset      => sdram_pll_reset_source_reset,     --    clk_reset.reset
			master_address       => jtag_master_master_address,       --       master.address
			master_readdata      => jtag_master_master_readdata,      --             .readdata
			master_read          => jtag_master_master_read,          --             .read
			master_write         => jtag_master_master_write,         --             .write
			master_writedata     => jtag_master_master_writedata,     --             .writedata
			master_waitrequest   => jtag_master_master_waitrequest,   --             .waitrequest
			master_readdatavalid => jtag_master_master_readdatavalid, --             .readdatavalid
			master_byteenable    => jtag_master_master_byteenable,    --             .byteenable
			master_reset_reset   => jtag_master_master_reset_reset    -- master_reset.reset
		);

	key : component AvalonMM_key
		port map (
			clk        => clk_clk,                                                     --                        clk.clk
			reset      => rst_controller_reset_out_reset,                              --                      reset.reset
			address    => mm_interconnect_0_key_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_key_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_key_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_key_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_key_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_key_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_key_avalon_parallel_port_slave_readdata,   --                           .readdata
			KEY        => pp_key_export                                                --         external_interface.export
		);

	led_g : component AvalonMM_led_g
		port map (
			clk        => clk_clk,                                                       --                        clk.clk
			reset      => rst_controller_reset_out_reset,                                --                      reset.reset
			address    => mm_interconnect_0_led_g_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_led_g_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_led_g_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_led_g_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_led_g_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_led_g_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_led_g_avalon_parallel_port_slave_readdata,   --                           .readdata
			LEDG       => pp_led_g_export                                                --         external_interface.export
		);

	led_r : component AvalonMM_led_r
		port map (
			clk        => clk_clk,                                                       --                        clk.clk
			reset      => rst_controller_reset_out_reset,                                --                      reset.reset
			address    => mm_interconnect_0_led_r_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_led_r_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_led_r_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_led_r_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_led_r_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_led_r_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_led_r_avalon_parallel_port_slave_readdata,   --                           .readdata
			LEDR       => pp_led_r_export                                                --         external_interface.export
		);

	mm_bridge : component altera_avalon_mm_bridge
		generic map (
			DATA_WIDTH        => 32,
			SYMBOL_WIDTH      => 8,
			HDL_ADDR_WIDTH    => 28,
			BURSTCOUNT_WIDTH  => 1,
			PIPELINE_COMMAND  => 0,
			PIPELINE_RESPONSE => 0
		)
		port map (
			clk              => sdram_pll_sys_clk_clk,              --   clk.clk
			reset            => rst_controller_001_reset_out_reset, -- reset.reset
			s0_waitrequest   => mm_bridge_s_waitrequest,            --    s0.waitrequest
			s0_readdata      => mm_bridge_s_readdata,               --      .readdata
			s0_readdatavalid => mm_bridge_s_readdatavalid,          --      .readdatavalid
			s0_burstcount    => mm_bridge_s_burstcount,             --      .burstcount
			s0_writedata     => mm_bridge_s_writedata,              --      .writedata
			s0_address       => mm_bridge_s_address,                --      .address
			s0_write         => mm_bridge_s_write,                  --      .write
			s0_read          => mm_bridge_s_read,                   --      .read
			s0_byteenable    => mm_bridge_s_byteenable,             --      .byteenable
			s0_debugaccess   => mm_bridge_s_debugaccess,            --      .debugaccess
			m0_waitrequest   => mm_bridge_m0_waitrequest,           --    m0.waitrequest
			m0_readdata      => mm_bridge_m0_readdata,              --      .readdata
			m0_readdatavalid => mm_bridge_m0_readdatavalid,         --      .readdatavalid
			m0_burstcount    => mm_bridge_m0_burstcount,            --      .burstcount
			m0_writedata     => mm_bridge_m0_writedata,             --      .writedata
			m0_address       => mm_bridge_m0_address,               --      .address
			m0_write         => mm_bridge_m0_write,                 --      .write
			m0_read          => mm_bridge_m0_read,                  --      .read
			m0_byteenable    => mm_bridge_m0_byteenable,            --      .byteenable
			m0_debugaccess   => mm_bridge_m0_debugaccess,           --      .debugaccess
			s0_response      => open,                               -- (terminated)
			m0_response      => "00"                                -- (terminated)
		);

	sdram_controller : component AvalonMM_sdram_controller
		port map (
			clk            => sdram_pll_sys_clk_clk,                                      --   clk.clk
			reset_n        => rst_controller_002_reset_out_reset_ports_inv,               -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_controller_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_controller_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_controller_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_controller_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_controller_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_controller_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_controller_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_controller_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                                 --  wire.export
			zs_ba          => sdram_ba,                                                   --      .export
			zs_cas_n       => sdram_cas_n,                                                --      .export
			zs_cke         => sdram_cke,                                                  --      .export
			zs_cs_n        => sdram_cs_n,                                                 --      .export
			zs_dq          => sdram_dq,                                                   --      .export
			zs_dqm         => sdram_dqm,                                                  --      .export
			zs_ras_n       => sdram_ras_n,                                                --      .export
			zs_we_n        => sdram_we_n                                                  --      .export
		);

	sdram_pll : component AvalonMM_sdram_pll
		port map (
			ref_clk_clk        => clk_clk,                        --      ref_clk.clk
			ref_reset_reset    => rst_controller_reset_out_reset, --    ref_reset.reset
			sys_clk_clk        => sdram_pll_sys_clk_clk,          --      sys_clk.clk
			sdram_clk_clk      => sdram_clk_clk,                  --    sdram_clk.clk
			reset_source_reset => sdram_pll_reset_source_reset    -- reset_source.reset
		);

	switch : component AvalonMM_switch
		port map (
			clk        => clk_clk,                                                        --                        clk.clk
			reset      => rst_controller_reset_out_reset,                                 --                      reset.reset
			address    => mm_interconnect_0_switch_avalon_parallel_port_slave_address,    -- avalon_parallel_port_slave.address
			byteenable => mm_interconnect_0_switch_avalon_parallel_port_slave_byteenable, --                           .byteenable
			chipselect => mm_interconnect_0_switch_avalon_parallel_port_slave_chipselect, --                           .chipselect
			read       => mm_interconnect_0_switch_avalon_parallel_port_slave_read,       --                           .read
			write      => mm_interconnect_0_switch_avalon_parallel_port_slave_write,      --                           .write
			writedata  => mm_interconnect_0_switch_avalon_parallel_port_slave_writedata,  --                           .writedata
			readdata   => mm_interconnect_0_switch_avalon_parallel_port_slave_readdata,   --                           .readdata
			SW         => pp_switch_export,                                               --         external_interface.export
			irq        => switch_int_irq                                                  --                  interrupt.irq
		);

	mm_interconnect_0 : component AvalonMM_mm_interconnect_0
		port map (
			clk_0_clk_clk                                      => clk_clk,                                                        --                                    clk_0_clk.clk
			sdram_pll_sys_clk_clk                              => sdram_pll_sys_clk_clk,                                          --                            sdram_pll_sys_clk.clk
			jtag_master_clk_reset_reset_bridge_in_reset_reset  => rst_controller_001_reset_out_reset,                             --  jtag_master_clk_reset_reset_bridge_in_reset.reset
			led_r_reset_reset_bridge_in_reset_reset            => rst_controller_reset_out_reset,                                 --            led_r_reset_reset_bridge_in_reset.reset
			mm_bridge_reset_reset_bridge_in_reset_reset        => rst_controller_001_reset_out_reset,                             --        mm_bridge_reset_reset_bridge_in_reset.reset
			sdram_controller_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                             -- sdram_controller_reset_reset_bridge_in_reset.reset
			jtag_master_master_address                         => jtag_master_master_address,                                     --                           jtag_master_master.address
			jtag_master_master_waitrequest                     => jtag_master_master_waitrequest,                                 --                                             .waitrequest
			jtag_master_master_byteenable                      => jtag_master_master_byteenable,                                  --                                             .byteenable
			jtag_master_master_read                            => jtag_master_master_read,                                        --                                             .read
			jtag_master_master_readdata                        => jtag_master_master_readdata,                                    --                                             .readdata
			jtag_master_master_readdatavalid                   => jtag_master_master_readdatavalid,                               --                                             .readdatavalid
			jtag_master_master_write                           => jtag_master_master_write,                                       --                                             .write
			jtag_master_master_writedata                       => jtag_master_master_writedata,                                   --                                             .writedata
			mm_bridge_m0_address                               => mm_bridge_m0_address,                                           --                                 mm_bridge_m0.address
			mm_bridge_m0_waitrequest                           => mm_bridge_m0_waitrequest,                                       --                                             .waitrequest
			mm_bridge_m0_burstcount                            => mm_bridge_m0_burstcount,                                        --                                             .burstcount
			mm_bridge_m0_byteenable                            => mm_bridge_m0_byteenable,                                        --                                             .byteenable
			mm_bridge_m0_read                                  => mm_bridge_m0_read,                                              --                                             .read
			mm_bridge_m0_readdata                              => mm_bridge_m0_readdata,                                          --                                             .readdata
			mm_bridge_m0_readdatavalid                         => mm_bridge_m0_readdatavalid,                                     --                                             .readdatavalid
			mm_bridge_m0_write                                 => mm_bridge_m0_write,                                             --                                             .write
			mm_bridge_m0_writedata                             => mm_bridge_m0_writedata,                                         --                                             .writedata
			mm_bridge_m0_debugaccess                           => mm_bridge_m0_debugaccess,                                       --                                             .debugaccess
			hex_03_avalon_parallel_port_slave_address          => mm_interconnect_0_hex_03_avalon_parallel_port_slave_address,    --            hex_03_avalon_parallel_port_slave.address
			hex_03_avalon_parallel_port_slave_write            => mm_interconnect_0_hex_03_avalon_parallel_port_slave_write,      --                                             .write
			hex_03_avalon_parallel_port_slave_read             => mm_interconnect_0_hex_03_avalon_parallel_port_slave_read,       --                                             .read
			hex_03_avalon_parallel_port_slave_readdata         => mm_interconnect_0_hex_03_avalon_parallel_port_slave_readdata,   --                                             .readdata
			hex_03_avalon_parallel_port_slave_writedata        => mm_interconnect_0_hex_03_avalon_parallel_port_slave_writedata,  --                                             .writedata
			hex_03_avalon_parallel_port_slave_byteenable       => mm_interconnect_0_hex_03_avalon_parallel_port_slave_byteenable, --                                             .byteenable
			hex_03_avalon_parallel_port_slave_chipselect       => mm_interconnect_0_hex_03_avalon_parallel_port_slave_chipselect, --                                             .chipselect
			hex_47_avalon_parallel_port_slave_address          => mm_interconnect_0_hex_47_avalon_parallel_port_slave_address,    --            hex_47_avalon_parallel_port_slave.address
			hex_47_avalon_parallel_port_slave_write            => mm_interconnect_0_hex_47_avalon_parallel_port_slave_write,      --                                             .write
			hex_47_avalon_parallel_port_slave_read             => mm_interconnect_0_hex_47_avalon_parallel_port_slave_read,       --                                             .read
			hex_47_avalon_parallel_port_slave_readdata         => mm_interconnect_0_hex_47_avalon_parallel_port_slave_readdata,   --                                             .readdata
			hex_47_avalon_parallel_port_slave_writedata        => mm_interconnect_0_hex_47_avalon_parallel_port_slave_writedata,  --                                             .writedata
			hex_47_avalon_parallel_port_slave_byteenable       => mm_interconnect_0_hex_47_avalon_parallel_port_slave_byteenable, --                                             .byteenable
			hex_47_avalon_parallel_port_slave_chipselect       => mm_interconnect_0_hex_47_avalon_parallel_port_slave_chipselect, --                                             .chipselect
			key_avalon_parallel_port_slave_address             => mm_interconnect_0_key_avalon_parallel_port_slave_address,       --               key_avalon_parallel_port_slave.address
			key_avalon_parallel_port_slave_write               => mm_interconnect_0_key_avalon_parallel_port_slave_write,         --                                             .write
			key_avalon_parallel_port_slave_read                => mm_interconnect_0_key_avalon_parallel_port_slave_read,          --                                             .read
			key_avalon_parallel_port_slave_readdata            => mm_interconnect_0_key_avalon_parallel_port_slave_readdata,      --                                             .readdata
			key_avalon_parallel_port_slave_writedata           => mm_interconnect_0_key_avalon_parallel_port_slave_writedata,     --                                             .writedata
			key_avalon_parallel_port_slave_byteenable          => mm_interconnect_0_key_avalon_parallel_port_slave_byteenable,    --                                             .byteenable
			key_avalon_parallel_port_slave_chipselect          => mm_interconnect_0_key_avalon_parallel_port_slave_chipselect,    --                                             .chipselect
			led_g_avalon_parallel_port_slave_address           => mm_interconnect_0_led_g_avalon_parallel_port_slave_address,     --             led_g_avalon_parallel_port_slave.address
			led_g_avalon_parallel_port_slave_write             => mm_interconnect_0_led_g_avalon_parallel_port_slave_write,       --                                             .write
			led_g_avalon_parallel_port_slave_read              => mm_interconnect_0_led_g_avalon_parallel_port_slave_read,        --                                             .read
			led_g_avalon_parallel_port_slave_readdata          => mm_interconnect_0_led_g_avalon_parallel_port_slave_readdata,    --                                             .readdata
			led_g_avalon_parallel_port_slave_writedata         => mm_interconnect_0_led_g_avalon_parallel_port_slave_writedata,   --                                             .writedata
			led_g_avalon_parallel_port_slave_byteenable        => mm_interconnect_0_led_g_avalon_parallel_port_slave_byteenable,  --                                             .byteenable
			led_g_avalon_parallel_port_slave_chipselect        => mm_interconnect_0_led_g_avalon_parallel_port_slave_chipselect,  --                                             .chipselect
			led_r_avalon_parallel_port_slave_address           => mm_interconnect_0_led_r_avalon_parallel_port_slave_address,     --             led_r_avalon_parallel_port_slave.address
			led_r_avalon_parallel_port_slave_write             => mm_interconnect_0_led_r_avalon_parallel_port_slave_write,       --                                             .write
			led_r_avalon_parallel_port_slave_read              => mm_interconnect_0_led_r_avalon_parallel_port_slave_read,        --                                             .read
			led_r_avalon_parallel_port_slave_readdata          => mm_interconnect_0_led_r_avalon_parallel_port_slave_readdata,    --                                             .readdata
			led_r_avalon_parallel_port_slave_writedata         => mm_interconnect_0_led_r_avalon_parallel_port_slave_writedata,   --                                             .writedata
			led_r_avalon_parallel_port_slave_byteenable        => mm_interconnect_0_led_r_avalon_parallel_port_slave_byteenable,  --                                             .byteenable
			led_r_avalon_parallel_port_slave_chipselect        => mm_interconnect_0_led_r_avalon_parallel_port_slave_chipselect,  --                                             .chipselect
			sdram_controller_s1_address                        => mm_interconnect_0_sdram_controller_s1_address,                  --                          sdram_controller_s1.address
			sdram_controller_s1_write                          => mm_interconnect_0_sdram_controller_s1_write,                    --                                             .write
			sdram_controller_s1_read                           => mm_interconnect_0_sdram_controller_s1_read,                     --                                             .read
			sdram_controller_s1_readdata                       => mm_interconnect_0_sdram_controller_s1_readdata,                 --                                             .readdata
			sdram_controller_s1_writedata                      => mm_interconnect_0_sdram_controller_s1_writedata,                --                                             .writedata
			sdram_controller_s1_byteenable                     => mm_interconnect_0_sdram_controller_s1_byteenable,               --                                             .byteenable
			sdram_controller_s1_readdatavalid                  => mm_interconnect_0_sdram_controller_s1_readdatavalid,            --                                             .readdatavalid
			sdram_controller_s1_waitrequest                    => mm_interconnect_0_sdram_controller_s1_waitrequest,              --                                             .waitrequest
			sdram_controller_s1_chipselect                     => mm_interconnect_0_sdram_controller_s1_chipselect,               --                                             .chipselect
			switch_avalon_parallel_port_slave_address          => mm_interconnect_0_switch_avalon_parallel_port_slave_address,    --            switch_avalon_parallel_port_slave.address
			switch_avalon_parallel_port_slave_write            => mm_interconnect_0_switch_avalon_parallel_port_slave_write,      --                                             .write
			switch_avalon_parallel_port_slave_read             => mm_interconnect_0_switch_avalon_parallel_port_slave_read,       --                                             .read
			switch_avalon_parallel_port_slave_readdata         => mm_interconnect_0_switch_avalon_parallel_port_slave_readdata,   --                                             .readdata
			switch_avalon_parallel_port_slave_writedata        => mm_interconnect_0_switch_avalon_parallel_port_slave_writedata,  --                                             .writedata
			switch_avalon_parallel_port_slave_byteenable       => mm_interconnect_0_switch_avalon_parallel_port_slave_byteenable, --                                             .byteenable
			switch_avalon_parallel_port_slave_chipselect       => mm_interconnect_0_switch_avalon_parallel_port_slave_chipselect  --                                             .chipselect
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => sdram_pll_reset_source_reset,       -- reset_in0.reset
			clk            => sdram_pll_sys_clk_clk,              --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => jtag_master_master_reset_reset,     -- reset_in0.reset
			clk            => sdram_pll_sys_clk_clk,              --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_sdram_controller_s1_read_ports_inv <= not mm_interconnect_0_sdram_controller_s1_read;

	mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_controller_s1_byteenable;

	mm_interconnect_0_sdram_controller_s1_write_ports_inv <= not mm_interconnect_0_sdram_controller_s1_write;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

end architecture rtl; -- of AvalonMM
