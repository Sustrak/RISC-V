-- AvalonMM.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity AvalonMM is
	port (
		clk_clk                   : in    std_logic                     := '0';             --           clk.clk
		mm_bridge_s_waitrequest   : out   std_logic;                                        --   mm_bridge_s.waitrequest
		mm_bridge_s_readdata      : out   std_logic_vector(31 downto 0);                    --              .readdata
		mm_bridge_s_readdatavalid : out   std_logic;                                        --              .readdatavalid
		mm_bridge_s_burstcount    : in    std_logic_vector(0 downto 0)  := (others => '0'); --              .burstcount
		mm_bridge_s_writedata     : in    std_logic_vector(31 downto 0) := (others => '0'); --              .writedata
		mm_bridge_s_address       : in    std_logic_vector(27 downto 0) := (others => '0'); --              .address
		mm_bridge_s_write         : in    std_logic                     := '0';             --              .write
		mm_bridge_s_read          : in    std_logic                     := '0';             --              .read
		mm_bridge_s_byteenable    : in    std_logic_vector(3 downto 0)  := (others => '0'); --              .byteenable
		mm_bridge_s_debugaccess   : in    std_logic                     := '0';             --              .debugaccess
		pp_key_export             : in    std_logic_vector(3 downto 0)  := (others => '0'); --        pp_key.export
		pp_key_int_irq            : out   std_logic;                                        --    pp_key_int.irq
		pp_led_g_export           : out   std_logic_vector(8 downto 0);                     --      pp_led_g.export
		pp_led_r_export           : out   std_logic_vector(17 downto 0);                    --      pp_led_r.export
		pp_sev_seg03_export       : out   std_logic_vector(31 downto 0);                    --  pp_sev_seg03.export
		pp_sev_seg47_export       : out   std_logic_vector(31 downto 0);                    --  pp_sev_seg47.export
		pp_switch_export          : in    std_logic_vector(17 downto 0) := (others => '0'); --     pp_switch.export
		pp_switch_int_irq         : out   std_logic;                                        -- pp_switch_int.irq
		ps2_CLK                   : inout std_logic                     := '0';             --           ps2.CLK
		ps2_DAT                   : inout std_logic                     := '0';             --              .DAT
		ps2_int_irq               : out   std_logic;                                        --       ps2_int.irq
		reset_reset_n             : in    std_logic                     := '0';             --         reset.reset_n
		sdram_addr                : out   std_logic_vector(12 downto 0);                    --         sdram.addr
		sdram_ba                  : out   std_logic_vector(1 downto 0);                     --              .ba
		sdram_cas_n               : out   std_logic;                                        --              .cas_n
		sdram_cke                 : out   std_logic;                                        --              .cke
		sdram_cs_n                : out   std_logic;                                        --              .cs_n
		sdram_dq                  : inout std_logic_vector(31 downto 0) := (others => '0'); --              .dq
		sdram_dqm                 : out   std_logic_vector(3 downto 0);                     --              .dqm
		sdram_ras_n               : out   std_logic;                                        --              .ras_n
		sdram_we_n                : out   std_logic;                                        --              .we_n
		sdram_clk_clk             : out   std_logic;                                        --     sdram_clk.clk
		sram_DQ                   : inout std_logic_vector(15 downto 0) := (others => '0'); --          sram.DQ
		sram_ADDR                 : out   std_logic_vector(19 downto 0);                    --              .ADDR
		sram_LB_N                 : out   std_logic;                                        --              .LB_N
		sram_UB_N                 : out   std_logic;                                        --              .UB_N
		sram_CE_N                 : out   std_logic;                                        --              .CE_N
		sram_OE_N                 : out   std_logic;                                        --              .OE_N
		sram_WE_N                 : out   std_logic;                                        --              .WE_N
		vga_CLK                   : out   std_logic;                                        --           vga.CLK
		vga_HS                    : out   std_logic;                                        --              .HS
		vga_VS                    : out   std_logic;                                        --              .VS
		vga_BLANK                 : out   std_logic;                                        --              .BLANK
		vga_SYNC                  : out   std_logic;                                        --              .SYNC
		vga_R                     : out   std_logic_vector(7 downto 0);                     --              .R
		vga_G                     : out   std_logic_vector(7 downto 0);                     --              .G
		vga_B                     : out   std_logic_vector(7 downto 0)                      --              .B
	);
end entity AvalonMM;

architecture rtl of AvalonMM is
	component AvalonMM_jtag_master is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component AvalonMM_jtag_master;

	component AvalonMM_key is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component AvalonMM_key;

	component AvalonMM_led_r is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(17 downto 0)                     -- export
		);
	end component AvalonMM_led_r;

	component AvalonMM_leg_g is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(8 downto 0)                      -- export
		);
	end component AvalonMM_leg_g;

	component altera_avalon_mm_bridge is
		generic (
			DATA_WIDTH        : integer := 32;
			SYMBOL_WIDTH      : integer := 8;
			HDL_ADDR_WIDTH    : integer := 10;
			BURSTCOUNT_WIDTH  : integer := 1;
			PIPELINE_COMMAND  : integer := 1;
			PIPELINE_RESPONSE : integer := 1
		);
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(27 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic;                                        -- debugaccess
			s0_response      : out std_logic_vector(1 downto 0);                     -- response
			m0_response      : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- response
		);
	end component altera_avalon_mm_bridge;

	component AvalonMM_ps2 is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic                     := 'X';             -- address
			chipselect  : in    std_logic                     := 'X';             -- chipselect
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			irq         : out   std_logic;                                        -- irq
			PS2_CLK     : inout std_logic                     := 'X';             -- export
			PS2_DAT     : inout std_logic                     := 'X'              -- export
		);
	end component AvalonMM_ps2;

	component AvalonMM_sdram_controller is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(31 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(31 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(3 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component AvalonMM_sdram_controller;

	component AvalonMM_sdram_pll is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component AvalonMM_sdram_pll;

	component AvalonMM_sev_seg03 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component AvalonMM_sev_seg03;

	component AvalonMM_sram_0 is
		port (
			clk           : in    std_logic                     := 'X';             -- clk
			reset         : in    std_logic                     := 'X';             -- reset
			SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			SRAM_ADDR     : out   std_logic_vector(19 downto 0);                    -- export
			SRAM_LB_N     : out   std_logic;                                        -- export
			SRAM_UB_N     : out   std_logic;                                        -- export
			SRAM_CE_N     : out   std_logic;                                        -- export
			SRAM_OE_N     : out   std_logic;                                        -- export
			SRAM_WE_N     : out   std_logic;                                        -- export
			address       : in    std_logic_vector(19 downto 0) := (others => 'X'); -- address
			byteenable    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			read          : in    std_logic                     := 'X';             -- read
			write         : in    std_logic                     := 'X';             -- write
			writedata     : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out   std_logic_vector(15 downto 0);                    -- readdata
			readdatavalid : out   std_logic                                         -- readdatavalid
		);
	end component AvalonMM_sram_0;

	component AvalonMM_switch is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(17 downto 0) := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component AvalonMM_switch;

	component AvalonMM_vga is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			data          : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			startofpacket : in  std_logic                     := 'X';             -- startofpacket
			endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			valid         : in  std_logic                     := 'X';             -- valid
			ready         : out std_logic;                                        -- ready
			VGA_CLK       : out std_logic;                                        -- export
			VGA_HS        : out std_logic;                                        -- export
			VGA_VS        : out std_logic;                                        -- export
			VGA_BLANK     : out std_logic;                                        -- export
			VGA_SYNC      : out std_logic;                                        -- export
			VGA_R         : out std_logic_vector(7 downto 0);                     -- export
			VGA_G         : out std_logic_vector(7 downto 0);                     -- export
			VGA_B         : out std_logic_vector(7 downto 0)                      -- export
		);
	end component AvalonMM_vga;

	component AvalonMM_vga_dma is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_arbiterlock   : out std_logic;                                        -- lock
			master_read          : out std_logic;                                        -- read
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_data          : out std_logic_vector(29 downto 0);                    -- data
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic                                         -- valid
		);
	end component AvalonMM_vga_dma;

	component AvalonMM_vga_pll is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			vga_clk_clk        : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component AvalonMM_vga_pll;

	component AvalonMM_video_dual_clock_buffer_0 is
		port (
			clk_stream_in            : in  std_logic                     := 'X';             -- clk
			reset_stream_in          : in  std_logic                     := 'X';             -- reset
			clk_stream_out           : in  std_logic                     := 'X';             -- clk
			reset_stream_out         : in  std_logic                     := 'X';             -- reset
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_data           : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component AvalonMM_video_dual_clock_buffer_0;

	component AvalonMM_mm_interconnect_0 is
		port (
			sdram_pll_sys_clk_clk                              : in  std_logic                     := 'X';             -- clk
			jtag_master_clk_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			sdram_controller_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			vga_dma_reset_reset_bridge_in_reset_reset          : in  std_logic                     := 'X';             -- reset
			jtag_master_master_address                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			jtag_master_master_waitrequest                     : out std_logic;                                        -- waitrequest
			jtag_master_master_byteenable                      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_master_master_read                            : in  std_logic                     := 'X';             -- read
			jtag_master_master_readdata                        : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_master_master_readdatavalid                   : out std_logic;                                        -- readdatavalid
			jtag_master_master_write                           : in  std_logic                     := 'X';             -- write
			jtag_master_master_writedata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			mm_bridge_m0_address                               : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			mm_bridge_m0_waitrequest                           : out std_logic;                                        -- waitrequest
			mm_bridge_m0_burstcount                            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			mm_bridge_m0_byteenable                            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			mm_bridge_m0_read                                  : in  std_logic                     := 'X';             -- read
			mm_bridge_m0_readdata                              : out std_logic_vector(31 downto 0);                    -- readdata
			mm_bridge_m0_readdatavalid                         : out std_logic;                                        -- readdatavalid
			mm_bridge_m0_write                                 : in  std_logic                     := 'X';             -- write
			mm_bridge_m0_writedata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			mm_bridge_m0_debugaccess                           : in  std_logic                     := 'X';             -- debugaccess
			vga_dma_avalon_dma_master_address                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			vga_dma_avalon_dma_master_waitrequest              : out std_logic;                                        -- waitrequest
			vga_dma_avalon_dma_master_read                     : in  std_logic                     := 'X';             -- read
			vga_dma_avalon_dma_master_readdata                 : out std_logic_vector(31 downto 0);                    -- readdata
			vga_dma_avalon_dma_master_readdatavalid            : out std_logic;                                        -- readdatavalid
			vga_dma_avalon_dma_master_lock                     : in  std_logic                     := 'X';             -- lock
			key_s1_address                                     : out std_logic_vector(1 downto 0);                     -- address
			key_s1_write                                       : out std_logic;                                        -- write
			key_s1_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			key_s1_writedata                                   : out std_logic_vector(31 downto 0);                    -- writedata
			key_s1_chipselect                                  : out std_logic;                                        -- chipselect
			led_r_s1_address                                   : out std_logic_vector(1 downto 0);                     -- address
			led_r_s1_write                                     : out std_logic;                                        -- write
			led_r_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_r_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			led_r_s1_chipselect                                : out std_logic;                                        -- chipselect
			leg_g_s1_address                                   : out std_logic_vector(1 downto 0);                     -- address
			leg_g_s1_write                                     : out std_logic;                                        -- write
			leg_g_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			leg_g_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			leg_g_s1_chipselect                                : out std_logic;                                        -- chipselect
			ps2_avalon_ps2_slave_address                       : out std_logic_vector(0 downto 0);                     -- address
			ps2_avalon_ps2_slave_write                         : out std_logic;                                        -- write
			ps2_avalon_ps2_slave_read                          : out std_logic;                                        -- read
			ps2_avalon_ps2_slave_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ps2_avalon_ps2_slave_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			ps2_avalon_ps2_slave_byteenable                    : out std_logic_vector(3 downto 0);                     -- byteenable
			ps2_avalon_ps2_slave_waitrequest                   : in  std_logic                     := 'X';             -- waitrequest
			ps2_avalon_ps2_slave_chipselect                    : out std_logic;                                        -- chipselect
			sdram_controller_s1_address                        : out std_logic_vector(24 downto 0);                    -- address
			sdram_controller_s1_write                          : out std_logic;                                        -- write
			sdram_controller_s1_read                           : out std_logic;                                        -- read
			sdram_controller_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sdram_controller_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			sdram_controller_s1_byteenable                     : out std_logic_vector(3 downto 0);                     -- byteenable
			sdram_controller_s1_readdatavalid                  : in  std_logic                     := 'X';             -- readdatavalid
			sdram_controller_s1_waitrequest                    : in  std_logic                     := 'X';             -- waitrequest
			sdram_controller_s1_chipselect                     : out std_logic;                                        -- chipselect
			sev_seg03_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			sev_seg03_s1_write                                 : out std_logic;                                        -- write
			sev_seg03_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sev_seg03_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			sev_seg03_s1_chipselect                            : out std_logic;                                        -- chipselect
			sev_seg47_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			sev_seg47_s1_write                                 : out std_logic;                                        -- write
			sev_seg47_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sev_seg47_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			sev_seg47_s1_chipselect                            : out std_logic;                                        -- chipselect
			sram_0_avalon_sram_slave_address                   : out std_logic_vector(19 downto 0);                    -- address
			sram_0_avalon_sram_slave_write                     : out std_logic;                                        -- write
			sram_0_avalon_sram_slave_read                      : out std_logic;                                        -- read
			sram_0_avalon_sram_slave_readdata                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sram_0_avalon_sram_slave_writedata                 : out std_logic_vector(15 downto 0);                    -- writedata
			sram_0_avalon_sram_slave_byteenable                : out std_logic_vector(1 downto 0);                     -- byteenable
			sram_0_avalon_sram_slave_readdatavalid             : in  std_logic                     := 'X';             -- readdatavalid
			switch_s1_address                                  : out std_logic_vector(1 downto 0);                     -- address
			switch_s1_write                                    : out std_logic;                                        -- write
			switch_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			switch_s1_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			switch_s1_chipselect                               : out std_logic;                                        -- chipselect
			vga_dma_avalon_dma_control_slave_address           : out std_logic_vector(1 downto 0);                     -- address
			vga_dma_avalon_dma_control_slave_write             : out std_logic;                                        -- write
			vga_dma_avalon_dma_control_slave_read              : out std_logic;                                        -- read
			vga_dma_avalon_dma_control_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			vga_dma_avalon_dma_control_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			vga_dma_avalon_dma_control_slave_byteenable        : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component AvalonMM_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal video_dual_clock_buffer_0_avalon_dc_buffer_source_valid         : std_logic;                     -- video_dual_clock_buffer_0:stream_out_valid -> vga:valid
	signal video_dual_clock_buffer_0_avalon_dc_buffer_source_data          : std_logic_vector(29 downto 0); -- video_dual_clock_buffer_0:stream_out_data -> vga:data
	signal video_dual_clock_buffer_0_avalon_dc_buffer_source_ready         : std_logic;                     -- vga:ready -> video_dual_clock_buffer_0:stream_out_ready
	signal video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket : std_logic;                     -- video_dual_clock_buffer_0:stream_out_startofpacket -> vga:startofpacket
	signal video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket   : std_logic;                     -- video_dual_clock_buffer_0:stream_out_endofpacket -> vga:endofpacket
	signal vga_dma_avalon_pixel_source_valid                               : std_logic;                     -- vga_dma:stream_valid -> video_dual_clock_buffer_0:stream_in_valid
	signal vga_dma_avalon_pixel_source_data                                : std_logic_vector(29 downto 0); -- vga_dma:stream_data -> video_dual_clock_buffer_0:stream_in_data
	signal vga_dma_avalon_pixel_source_ready                               : std_logic;                     -- video_dual_clock_buffer_0:stream_in_ready -> vga_dma:stream_ready
	signal vga_dma_avalon_pixel_source_startofpacket                       : std_logic;                     -- vga_dma:stream_startofpacket -> video_dual_clock_buffer_0:stream_in_startofpacket
	signal vga_dma_avalon_pixel_source_endofpacket                         : std_logic;                     -- vga_dma:stream_endofpacket -> video_dual_clock_buffer_0:stream_in_endofpacket
	signal sdram_pll_sys_clk_clk                                           : std_logic;                     -- sdram_pll:sys_clk_clk -> [jtag_master:clk_clk, key:clk, led_r:clk, leg_g:clk, mm_bridge:clk, mm_interconnect_0:sdram_pll_sys_clk_clk, ps2:clk, rst_controller:clk, rst_controller_001:clk, sdram_controller:clk, sev_seg03:clk, sev_seg47:clk, sram_0:clk, switch:clk, vga_dma:clk, vga_pll:ref_clk_clk, video_dual_clock_buffer_0:clk_stream_in]
	signal vga_pll_vga_clk_clk                                             : std_logic;                     -- vga_pll:vga_clk_clk -> [rst_controller_003:clk, vga:clk, video_dual_clock_buffer_0:clk_stream_out]
	signal sdram_pll_reset_source_reset                                    : std_logic;                     -- sdram_pll:reset_source_reset -> [jtag_master:clk_reset_reset, rst_controller:reset_in0]
	signal vga_dma_avalon_dma_master_waitrequest                           : std_logic;                     -- mm_interconnect_0:vga_dma_avalon_dma_master_waitrequest -> vga_dma:master_waitrequest
	signal vga_dma_avalon_dma_master_readdata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:vga_dma_avalon_dma_master_readdata -> vga_dma:master_readdata
	signal vga_dma_avalon_dma_master_address                               : std_logic_vector(31 downto 0); -- vga_dma:master_address -> mm_interconnect_0:vga_dma_avalon_dma_master_address
	signal vga_dma_avalon_dma_master_read                                  : std_logic;                     -- vga_dma:master_read -> mm_interconnect_0:vga_dma_avalon_dma_master_read
	signal vga_dma_avalon_dma_master_readdatavalid                         : std_logic;                     -- mm_interconnect_0:vga_dma_avalon_dma_master_readdatavalid -> vga_dma:master_readdatavalid
	signal vga_dma_avalon_dma_master_lock                                  : std_logic;                     -- vga_dma:master_arbiterlock -> mm_interconnect_0:vga_dma_avalon_dma_master_lock
	signal mm_bridge_m0_waitrequest                                        : std_logic;                     -- mm_interconnect_0:mm_bridge_m0_waitrequest -> mm_bridge:m0_waitrequest
	signal mm_bridge_m0_readdata                                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:mm_bridge_m0_readdata -> mm_bridge:m0_readdata
	signal mm_bridge_m0_debugaccess                                        : std_logic;                     -- mm_bridge:m0_debugaccess -> mm_interconnect_0:mm_bridge_m0_debugaccess
	signal mm_bridge_m0_address                                            : std_logic_vector(27 downto 0); -- mm_bridge:m0_address -> mm_interconnect_0:mm_bridge_m0_address
	signal mm_bridge_m0_read                                               : std_logic;                     -- mm_bridge:m0_read -> mm_interconnect_0:mm_bridge_m0_read
	signal mm_bridge_m0_byteenable                                         : std_logic_vector(3 downto 0);  -- mm_bridge:m0_byteenable -> mm_interconnect_0:mm_bridge_m0_byteenable
	signal mm_bridge_m0_readdatavalid                                      : std_logic;                     -- mm_interconnect_0:mm_bridge_m0_readdatavalid -> mm_bridge:m0_readdatavalid
	signal mm_bridge_m0_writedata                                          : std_logic_vector(31 downto 0); -- mm_bridge:m0_writedata -> mm_interconnect_0:mm_bridge_m0_writedata
	signal mm_bridge_m0_write                                              : std_logic;                     -- mm_bridge:m0_write -> mm_interconnect_0:mm_bridge_m0_write
	signal mm_bridge_m0_burstcount                                         : std_logic_vector(0 downto 0);  -- mm_bridge:m0_burstcount -> mm_interconnect_0:mm_bridge_m0_burstcount
	signal jtag_master_master_readdata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_master_master_readdata -> jtag_master:master_readdata
	signal jtag_master_master_waitrequest                                  : std_logic;                     -- mm_interconnect_0:jtag_master_master_waitrequest -> jtag_master:master_waitrequest
	signal jtag_master_master_address                                      : std_logic_vector(31 downto 0); -- jtag_master:master_address -> mm_interconnect_0:jtag_master_master_address
	signal jtag_master_master_read                                         : std_logic;                     -- jtag_master:master_read -> mm_interconnect_0:jtag_master_master_read
	signal jtag_master_master_byteenable                                   : std_logic_vector(3 downto 0);  -- jtag_master:master_byteenable -> mm_interconnect_0:jtag_master_master_byteenable
	signal jtag_master_master_readdatavalid                                : std_logic;                     -- mm_interconnect_0:jtag_master_master_readdatavalid -> jtag_master:master_readdatavalid
	signal jtag_master_master_write                                        : std_logic;                     -- jtag_master:master_write -> mm_interconnect_0:jtag_master_master_write
	signal jtag_master_master_writedata                                    : std_logic_vector(31 downto 0); -- jtag_master:master_writedata -> mm_interconnect_0:jtag_master_master_writedata
	signal mm_interconnect_0_sram_0_avalon_sram_slave_readdata             : std_logic_vector(15 downto 0); -- sram_0:readdata -> mm_interconnect_0:sram_0_avalon_sram_slave_readdata
	signal mm_interconnect_0_sram_0_avalon_sram_slave_address              : std_logic_vector(19 downto 0); -- mm_interconnect_0:sram_0_avalon_sram_slave_address -> sram_0:address
	signal mm_interconnect_0_sram_0_avalon_sram_slave_read                 : std_logic;                     -- mm_interconnect_0:sram_0_avalon_sram_slave_read -> sram_0:read
	signal mm_interconnect_0_sram_0_avalon_sram_slave_byteenable           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sram_0_avalon_sram_slave_byteenable -> sram_0:byteenable
	signal mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid        : std_logic;                     -- sram_0:readdatavalid -> mm_interconnect_0:sram_0_avalon_sram_slave_readdatavalid
	signal mm_interconnect_0_sram_0_avalon_sram_slave_write                : std_logic;                     -- mm_interconnect_0:sram_0_avalon_sram_slave_write -> sram_0:write
	signal mm_interconnect_0_sram_0_avalon_sram_slave_writedata            : std_logic_vector(15 downto 0); -- mm_interconnect_0:sram_0_avalon_sram_slave_writedata -> sram_0:writedata
	signal mm_interconnect_0_vga_dma_avalon_dma_control_slave_readdata     : std_logic_vector(31 downto 0); -- vga_dma:slave_readdata -> mm_interconnect_0:vga_dma_avalon_dma_control_slave_readdata
	signal mm_interconnect_0_vga_dma_avalon_dma_control_slave_address      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:vga_dma_avalon_dma_control_slave_address -> vga_dma:slave_address
	signal mm_interconnect_0_vga_dma_avalon_dma_control_slave_read         : std_logic;                     -- mm_interconnect_0:vga_dma_avalon_dma_control_slave_read -> vga_dma:slave_read
	signal mm_interconnect_0_vga_dma_avalon_dma_control_slave_byteenable   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:vga_dma_avalon_dma_control_slave_byteenable -> vga_dma:slave_byteenable
	signal mm_interconnect_0_vga_dma_avalon_dma_control_slave_write        : std_logic;                     -- mm_interconnect_0:vga_dma_avalon_dma_control_slave_write -> vga_dma:slave_write
	signal mm_interconnect_0_vga_dma_avalon_dma_control_slave_writedata    : std_logic_vector(31 downto 0); -- mm_interconnect_0:vga_dma_avalon_dma_control_slave_writedata -> vga_dma:slave_writedata
	signal mm_interconnect_0_ps2_avalon_ps2_slave_chipselect               : std_logic;                     -- mm_interconnect_0:ps2_avalon_ps2_slave_chipselect -> ps2:chipselect
	signal mm_interconnect_0_ps2_avalon_ps2_slave_readdata                 : std_logic_vector(31 downto 0); -- ps2:readdata -> mm_interconnect_0:ps2_avalon_ps2_slave_readdata
	signal mm_interconnect_0_ps2_avalon_ps2_slave_waitrequest              : std_logic;                     -- ps2:waitrequest -> mm_interconnect_0:ps2_avalon_ps2_slave_waitrequest
	signal mm_interconnect_0_ps2_avalon_ps2_slave_address                  : std_logic_vector(0 downto 0);  -- mm_interconnect_0:ps2_avalon_ps2_slave_address -> ps2:address
	signal mm_interconnect_0_ps2_avalon_ps2_slave_read                     : std_logic;                     -- mm_interconnect_0:ps2_avalon_ps2_slave_read -> ps2:read
	signal mm_interconnect_0_ps2_avalon_ps2_slave_byteenable               : std_logic_vector(3 downto 0);  -- mm_interconnect_0:ps2_avalon_ps2_slave_byteenable -> ps2:byteenable
	signal mm_interconnect_0_ps2_avalon_ps2_slave_write                    : std_logic;                     -- mm_interconnect_0:ps2_avalon_ps2_slave_write -> ps2:write
	signal mm_interconnect_0_ps2_avalon_ps2_slave_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:ps2_avalon_ps2_slave_writedata -> ps2:writedata
	signal mm_interconnect_0_sdram_controller_s1_chipselect                : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	signal mm_interconnect_0_sdram_controller_s1_readdata                  : std_logic_vector(31 downto 0); -- sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	signal mm_interconnect_0_sdram_controller_s1_waitrequest               : std_logic;                     -- sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	signal mm_interconnect_0_sdram_controller_s1_address                   : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	signal mm_interconnect_0_sdram_controller_s1_read                      : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_read -> mm_interconnect_0_sdram_controller_s1_read:in
	signal mm_interconnect_0_sdram_controller_s1_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:sdram_controller_s1_byteenable -> mm_interconnect_0_sdram_controller_s1_byteenable:in
	signal mm_interconnect_0_sdram_controller_s1_readdatavalid             : std_logic;                     -- sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	signal mm_interconnect_0_sdram_controller_s1_write                     : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_write -> mm_interconnect_0_sdram_controller_s1_write:in
	signal mm_interconnect_0_sdram_controller_s1_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	signal mm_interconnect_0_leg_g_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:leg_g_s1_chipselect -> leg_g:chipselect
	signal mm_interconnect_0_leg_g_s1_readdata                             : std_logic_vector(31 downto 0); -- leg_g:readdata -> mm_interconnect_0:leg_g_s1_readdata
	signal mm_interconnect_0_leg_g_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:leg_g_s1_address -> leg_g:address
	signal mm_interconnect_0_leg_g_s1_write                                : std_logic;                     -- mm_interconnect_0:leg_g_s1_write -> mm_interconnect_0_leg_g_s1_write:in
	signal mm_interconnect_0_leg_g_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:leg_g_s1_writedata -> leg_g:writedata
	signal mm_interconnect_0_switch_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:switch_s1_chipselect -> switch:chipselect
	signal mm_interconnect_0_switch_s1_readdata                            : std_logic_vector(31 downto 0); -- switch:readdata -> mm_interconnect_0:switch_s1_readdata
	signal mm_interconnect_0_switch_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switch_s1_address -> switch:address
	signal mm_interconnect_0_switch_s1_write                               : std_logic;                     -- mm_interconnect_0:switch_s1_write -> mm_interconnect_0_switch_s1_write:in
	signal mm_interconnect_0_switch_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:switch_s1_writedata -> switch:writedata
	signal mm_interconnect_0_key_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:key_s1_chipselect -> key:chipselect
	signal mm_interconnect_0_key_s1_readdata                               : std_logic_vector(31 downto 0); -- key:readdata -> mm_interconnect_0:key_s1_readdata
	signal mm_interconnect_0_key_s1_address                                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:key_s1_address -> key:address
	signal mm_interconnect_0_key_s1_write                                  : std_logic;                     -- mm_interconnect_0:key_s1_write -> mm_interconnect_0_key_s1_write:in
	signal mm_interconnect_0_key_s1_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:key_s1_writedata -> key:writedata
	signal mm_interconnect_0_led_r_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:led_r_s1_chipselect -> led_r:chipselect
	signal mm_interconnect_0_led_r_s1_readdata                             : std_logic_vector(31 downto 0); -- led_r:readdata -> mm_interconnect_0:led_r_s1_readdata
	signal mm_interconnect_0_led_r_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_r_s1_address -> led_r:address
	signal mm_interconnect_0_led_r_s1_write                                : std_logic;                     -- mm_interconnect_0:led_r_s1_write -> mm_interconnect_0_led_r_s1_write:in
	signal mm_interconnect_0_led_r_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_r_s1_writedata -> led_r:writedata
	signal mm_interconnect_0_sev_seg03_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:sev_seg03_s1_chipselect -> sev_seg03:chipselect
	signal mm_interconnect_0_sev_seg03_s1_readdata                         : std_logic_vector(31 downto 0); -- sev_seg03:readdata -> mm_interconnect_0:sev_seg03_s1_readdata
	signal mm_interconnect_0_sev_seg03_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sev_seg03_s1_address -> sev_seg03:address
	signal mm_interconnect_0_sev_seg03_s1_write                            : std_logic;                     -- mm_interconnect_0:sev_seg03_s1_write -> mm_interconnect_0_sev_seg03_s1_write:in
	signal mm_interconnect_0_sev_seg03_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:sev_seg03_s1_writedata -> sev_seg03:writedata
	signal mm_interconnect_0_sev_seg47_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:sev_seg47_s1_chipselect -> sev_seg47:chipselect
	signal mm_interconnect_0_sev_seg47_s1_readdata                         : std_logic_vector(31 downto 0); -- sev_seg47:readdata -> mm_interconnect_0:sev_seg47_s1_readdata
	signal mm_interconnect_0_sev_seg47_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sev_seg47_s1_address -> sev_seg47:address
	signal mm_interconnect_0_sev_seg47_s1_write                            : std_logic;                     -- mm_interconnect_0:sev_seg47_s1_write -> mm_interconnect_0_sev_seg47_s1_write:in
	signal mm_interconnect_0_sev_seg47_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:sev_seg47_s1_writedata -> sev_seg47:writedata
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [mm_bridge:reset, mm_interconnect_0:jtag_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:vga_dma_reset_reset_bridge_in_reset_reset, ps2:reset, rst_controller_reset_out_reset:in, sram_0:reset, vga_dma:reset, vga_pll:ref_reset_reset, video_dual_clock_buffer_0:reset_stream_in]
	signal rst_controller_001_reset_out_reset                              : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:sdram_controller_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal jtag_master_master_reset_reset                                  : std_logic;                     -- jtag_master:master_reset_reset -> rst_controller_001:reset_in0
	signal rst_controller_002_reset_out_reset                              : std_logic;                     -- rst_controller_002:reset_out -> sdram_pll:ref_reset_reset
	signal rst_controller_003_reset_out_reset                              : std_logic;                     -- rst_controller_003:reset_out -> [vga:reset, video_dual_clock_buffer_0:reset_stream_out]
	signal vga_pll_reset_source_reset                                      : std_logic;                     -- vga_pll:reset_source_reset -> rst_controller_003:reset_in0
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> rst_controller_002:reset_in0
	signal mm_interconnect_0_sdram_controller_s1_read_ports_inv            : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_read:inv -> sdram_controller:az_rd_n
	signal mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv      : std_logic_vector(3 downto 0);  -- mm_interconnect_0_sdram_controller_s1_byteenable:inv -> sdram_controller:az_be_n
	signal mm_interconnect_0_sdram_controller_s1_write_ports_inv           : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_write:inv -> sdram_controller:az_wr_n
	signal mm_interconnect_0_leg_g_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_leg_g_s1_write:inv -> leg_g:write_n
	signal mm_interconnect_0_switch_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_switch_s1_write:inv -> switch:write_n
	signal mm_interconnect_0_key_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_key_s1_write:inv -> key:write_n
	signal mm_interconnect_0_led_r_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_led_r_s1_write:inv -> led_r:write_n
	signal mm_interconnect_0_sev_seg03_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_sev_seg03_s1_write:inv -> sev_seg03:write_n
	signal mm_interconnect_0_sev_seg47_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_sev_seg47_s1_write:inv -> sev_seg47:write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [key:reset_n, led_r:reset_n, leg_g:reset_n, sev_seg03:reset_n, sev_seg47:reset_n, switch:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                    : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> sdram_controller:reset_n

begin

	jtag_master : component AvalonMM_jtag_master
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => sdram_pll_sys_clk_clk,            --          clk.clk
			clk_reset_reset      => sdram_pll_reset_source_reset,     --    clk_reset.reset
			master_address       => jtag_master_master_address,       --       master.address
			master_readdata      => jtag_master_master_readdata,      --             .readdata
			master_read          => jtag_master_master_read,          --             .read
			master_write         => jtag_master_master_write,         --             .write
			master_writedata     => jtag_master_master_writedata,     --             .writedata
			master_waitrequest   => jtag_master_master_waitrequest,   --             .waitrequest
			master_readdatavalid => jtag_master_master_readdatavalid, --             .readdatavalid
			master_byteenable    => jtag_master_master_byteenable,    --             .byteenable
			master_reset_reset   => jtag_master_master_reset_reset    -- master_reset.reset
		);

	key : component AvalonMM_key
		port map (
			clk        => sdram_pll_sys_clk_clk,                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_key_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_key_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_key_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_key_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_key_s1_readdata,        --                    .readdata
			in_port    => pp_key_export,                            -- external_connection.export
			irq        => pp_key_int_irq                            --                 irq.irq
		);

	led_r : component AvalonMM_led_r
		port map (
			clk        => sdram_pll_sys_clk_clk,                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_led_r_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_r_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_r_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_r_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_r_s1_readdata,        --                    .readdata
			out_port   => pp_led_r_export                             -- external_connection.export
		);

	leg_g : component AvalonMM_leg_g
		port map (
			clk        => sdram_pll_sys_clk_clk,                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_leg_g_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_leg_g_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_leg_g_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_leg_g_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_leg_g_s1_readdata,        --                    .readdata
			out_port   => pp_led_g_export                             -- external_connection.export
		);

	mm_bridge : component altera_avalon_mm_bridge
		generic map (
			DATA_WIDTH        => 32,
			SYMBOL_WIDTH      => 8,
			HDL_ADDR_WIDTH    => 28,
			BURSTCOUNT_WIDTH  => 1,
			PIPELINE_COMMAND  => 0,
			PIPELINE_RESPONSE => 0
		)
		port map (
			clk              => sdram_pll_sys_clk_clk,          --   clk.clk
			reset            => rst_controller_reset_out_reset, -- reset.reset
			s0_waitrequest   => mm_bridge_s_waitrequest,        --    s0.waitrequest
			s0_readdata      => mm_bridge_s_readdata,           --      .readdata
			s0_readdatavalid => mm_bridge_s_readdatavalid,      --      .readdatavalid
			s0_burstcount    => mm_bridge_s_burstcount,         --      .burstcount
			s0_writedata     => mm_bridge_s_writedata,          --      .writedata
			s0_address       => mm_bridge_s_address,            --      .address
			s0_write         => mm_bridge_s_write,              --      .write
			s0_read          => mm_bridge_s_read,               --      .read
			s0_byteenable    => mm_bridge_s_byteenable,         --      .byteenable
			s0_debugaccess   => mm_bridge_s_debugaccess,        --      .debugaccess
			m0_waitrequest   => mm_bridge_m0_waitrequest,       --    m0.waitrequest
			m0_readdata      => mm_bridge_m0_readdata,          --      .readdata
			m0_readdatavalid => mm_bridge_m0_readdatavalid,     --      .readdatavalid
			m0_burstcount    => mm_bridge_m0_burstcount,        --      .burstcount
			m0_writedata     => mm_bridge_m0_writedata,         --      .writedata
			m0_address       => mm_bridge_m0_address,           --      .address
			m0_write         => mm_bridge_m0_write,             --      .write
			m0_read          => mm_bridge_m0_read,              --      .read
			m0_byteenable    => mm_bridge_m0_byteenable,        --      .byteenable
			m0_debugaccess   => mm_bridge_m0_debugaccess,       --      .debugaccess
			s0_response      => open,                           -- (terminated)
			m0_response      => "00"                            -- (terminated)
		);

	ps2 : component AvalonMM_ps2
		port map (
			clk         => sdram_pll_sys_clk_clk,                              --                clk.clk
			reset       => rst_controller_reset_out_reset,                     --              reset.reset
			address     => mm_interconnect_0_ps2_avalon_ps2_slave_address(0),  --   avalon_ps2_slave.address
			chipselect  => mm_interconnect_0_ps2_avalon_ps2_slave_chipselect,  --                   .chipselect
			byteenable  => mm_interconnect_0_ps2_avalon_ps2_slave_byteenable,  --                   .byteenable
			read        => mm_interconnect_0_ps2_avalon_ps2_slave_read,        --                   .read
			write       => mm_interconnect_0_ps2_avalon_ps2_slave_write,       --                   .write
			writedata   => mm_interconnect_0_ps2_avalon_ps2_slave_writedata,   --                   .writedata
			readdata    => mm_interconnect_0_ps2_avalon_ps2_slave_readdata,    --                   .readdata
			waitrequest => mm_interconnect_0_ps2_avalon_ps2_slave_waitrequest, --                   .waitrequest
			irq         => ps2_int_irq,                                        --          interrupt.irq
			PS2_CLK     => ps2_CLK,                                            -- external_interface.export
			PS2_DAT     => ps2_DAT                                             --                   .export
		);

	sdram_controller : component AvalonMM_sdram_controller
		port map (
			clk            => sdram_pll_sys_clk_clk,                                      --   clk.clk
			reset_n        => rst_controller_001_reset_out_reset_ports_inv,               -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_controller_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_controller_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_controller_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_controller_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_controller_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_controller_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_controller_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_controller_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                                 --  wire.export
			zs_ba          => sdram_ba,                                                   --      .export
			zs_cas_n       => sdram_cas_n,                                                --      .export
			zs_cke         => sdram_cke,                                                  --      .export
			zs_cs_n        => sdram_cs_n,                                                 --      .export
			zs_dq          => sdram_dq,                                                   --      .export
			zs_dqm         => sdram_dqm,                                                  --      .export
			zs_ras_n       => sdram_ras_n,                                                --      .export
			zs_we_n        => sdram_we_n                                                  --      .export
		);

	sdram_pll : component AvalonMM_sdram_pll
		port map (
			ref_clk_clk        => clk_clk,                            --      ref_clk.clk
			ref_reset_reset    => rst_controller_002_reset_out_reset, --    ref_reset.reset
			sys_clk_clk        => sdram_pll_sys_clk_clk,              --      sys_clk.clk
			sdram_clk_clk      => sdram_clk_clk,                      --    sdram_clk.clk
			reset_source_reset => sdram_pll_reset_source_reset        -- reset_source.reset
		);

	sev_seg03 : component AvalonMM_sev_seg03
		port map (
			clk        => sdram_pll_sys_clk_clk,                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_sev_seg03_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_sev_seg03_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_sev_seg03_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_sev_seg03_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_sev_seg03_s1_readdata,        --                    .readdata
			out_port   => pp_sev_seg03_export                             -- external_connection.export
		);

	sev_seg47 : component AvalonMM_sev_seg03
		port map (
			clk        => sdram_pll_sys_clk_clk,                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_sev_seg47_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_sev_seg47_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_sev_seg47_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_sev_seg47_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_sev_seg47_s1_readdata,        --                    .readdata
			out_port   => pp_sev_seg47_export                             -- external_connection.export
		);

	sram_0 : component AvalonMM_sram_0
		port map (
			clk           => sdram_pll_sys_clk_clk,                                    --                clk.clk
			reset         => rst_controller_reset_out_reset,                           --              reset.reset
			SRAM_DQ       => sram_DQ,                                                  -- external_interface.export
			SRAM_ADDR     => sram_ADDR,                                                --                   .export
			SRAM_LB_N     => sram_LB_N,                                                --                   .export
			SRAM_UB_N     => sram_UB_N,                                                --                   .export
			SRAM_CE_N     => sram_CE_N,                                                --                   .export
			SRAM_OE_N     => sram_OE_N,                                                --                   .export
			SRAM_WE_N     => sram_WE_N,                                                --                   .export
			address       => mm_interconnect_0_sram_0_avalon_sram_slave_address,       --  avalon_sram_slave.address
			byteenable    => mm_interconnect_0_sram_0_avalon_sram_slave_byteenable,    --                   .byteenable
			read          => mm_interconnect_0_sram_0_avalon_sram_slave_read,          --                   .read
			write         => mm_interconnect_0_sram_0_avalon_sram_slave_write,         --                   .write
			writedata     => mm_interconnect_0_sram_0_avalon_sram_slave_writedata,     --                   .writedata
			readdata      => mm_interconnect_0_sram_0_avalon_sram_slave_readdata,      --                   .readdata
			readdatavalid => mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid  --                   .readdatavalid
		);

	switch : component AvalonMM_switch
		port map (
			clk        => sdram_pll_sys_clk_clk,                       --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_switch_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_switch_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_switch_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_switch_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_switch_s1_readdata,        --                    .readdata
			in_port    => pp_switch_export,                            -- external_connection.export
			irq        => pp_switch_int_irq                            --                 irq.irq
		);

	vga : component AvalonMM_vga
		port map (
			clk           => vga_pll_vga_clk_clk,                                             --                clk.clk
			reset         => rst_controller_003_reset_out_reset,                              --              reset.reset
			data          => video_dual_clock_buffer_0_avalon_dc_buffer_source_data,          --    avalon_vga_sink.data
			startofpacket => video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket, --                   .startofpacket
			endofpacket   => video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket,   --                   .endofpacket
			valid         => video_dual_clock_buffer_0_avalon_dc_buffer_source_valid,         --                   .valid
			ready         => video_dual_clock_buffer_0_avalon_dc_buffer_source_ready,         --                   .ready
			VGA_CLK       => vga_CLK,                                                         -- external_interface.export
			VGA_HS        => vga_HS,                                                          --                   .export
			VGA_VS        => vga_VS,                                                          --                   .export
			VGA_BLANK     => vga_BLANK,                                                       --                   .export
			VGA_SYNC      => vga_SYNC,                                                        --                   .export
			VGA_R         => vga_R,                                                           --                   .export
			VGA_G         => vga_G,                                                           --                   .export
			VGA_B         => vga_B                                                            --                   .export
		);

	vga_dma : component AvalonMM_vga_dma
		port map (
			clk                  => sdram_pll_sys_clk_clk,                                         --                      clk.clk
			reset                => rst_controller_reset_out_reset,                                --                    reset.reset
			master_address       => vga_dma_avalon_dma_master_address,                             --        avalon_dma_master.address
			master_waitrequest   => vga_dma_avalon_dma_master_waitrequest,                         --                         .waitrequest
			master_arbiterlock   => vga_dma_avalon_dma_master_lock,                                --                         .lock
			master_read          => vga_dma_avalon_dma_master_read,                                --                         .read
			master_readdata      => vga_dma_avalon_dma_master_readdata,                            --                         .readdata
			master_readdatavalid => vga_dma_avalon_dma_master_readdatavalid,                       --                         .readdatavalid
			slave_address        => mm_interconnect_0_vga_dma_avalon_dma_control_slave_address,    -- avalon_dma_control_slave.address
			slave_byteenable     => mm_interconnect_0_vga_dma_avalon_dma_control_slave_byteenable, --                         .byteenable
			slave_read           => mm_interconnect_0_vga_dma_avalon_dma_control_slave_read,       --                         .read
			slave_write          => mm_interconnect_0_vga_dma_avalon_dma_control_slave_write,      --                         .write
			slave_writedata      => mm_interconnect_0_vga_dma_avalon_dma_control_slave_writedata,  --                         .writedata
			slave_readdata       => mm_interconnect_0_vga_dma_avalon_dma_control_slave_readdata,   --                         .readdata
			stream_ready         => vga_dma_avalon_pixel_source_ready,                             --      avalon_pixel_source.ready
			stream_data          => vga_dma_avalon_pixel_source_data,                              --                         .data
			stream_startofpacket => vga_dma_avalon_pixel_source_startofpacket,                     --                         .startofpacket
			stream_endofpacket   => vga_dma_avalon_pixel_source_endofpacket,                       --                         .endofpacket
			stream_valid         => vga_dma_avalon_pixel_source_valid                              --                         .valid
		);

	vga_pll : component AvalonMM_vga_pll
		port map (
			ref_clk_clk        => sdram_pll_sys_clk_clk,          --      ref_clk.clk
			ref_reset_reset    => rst_controller_reset_out_reset, --    ref_reset.reset
			vga_clk_clk        => vga_pll_vga_clk_clk,            --      vga_clk.clk
			reset_source_reset => vga_pll_reset_source_reset      -- reset_source.reset
		);

	video_dual_clock_buffer_0 : component AvalonMM_video_dual_clock_buffer_0
		port map (
			clk_stream_in            => sdram_pll_sys_clk_clk,                                           --         clock_stream_in.clk
			reset_stream_in          => rst_controller_reset_out_reset,                                  --         reset_stream_in.reset
			clk_stream_out           => vga_pll_vga_clk_clk,                                             --        clock_stream_out.clk
			reset_stream_out         => rst_controller_003_reset_out_reset,                              --        reset_stream_out.reset
			stream_in_ready          => vga_dma_avalon_pixel_source_ready,                               --   avalon_dc_buffer_sink.ready
			stream_in_startofpacket  => vga_dma_avalon_pixel_source_startofpacket,                       --                        .startofpacket
			stream_in_endofpacket    => vga_dma_avalon_pixel_source_endofpacket,                         --                        .endofpacket
			stream_in_valid          => vga_dma_avalon_pixel_source_valid,                               --                        .valid
			stream_in_data           => vga_dma_avalon_pixel_source_data,                                --                        .data
			stream_out_ready         => video_dual_clock_buffer_0_avalon_dc_buffer_source_ready,         -- avalon_dc_buffer_source.ready
			stream_out_startofpacket => video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket, --                        .startofpacket
			stream_out_endofpacket   => video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket,   --                        .endofpacket
			stream_out_valid         => video_dual_clock_buffer_0_avalon_dc_buffer_source_valid,         --                        .valid
			stream_out_data          => video_dual_clock_buffer_0_avalon_dc_buffer_source_data           --                        .data
		);

	mm_interconnect_0 : component AvalonMM_mm_interconnect_0
		port map (
			sdram_pll_sys_clk_clk                              => sdram_pll_sys_clk_clk,                                         --                            sdram_pll_sys_clk.clk
			jtag_master_clk_reset_reset_bridge_in_reset_reset  => rst_controller_reset_out_reset,                                --  jtag_master_clk_reset_reset_bridge_in_reset.reset
			sdram_controller_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                            -- sdram_controller_reset_reset_bridge_in_reset.reset
			vga_dma_reset_reset_bridge_in_reset_reset          => rst_controller_reset_out_reset,                                --          vga_dma_reset_reset_bridge_in_reset.reset
			jtag_master_master_address                         => jtag_master_master_address,                                    --                           jtag_master_master.address
			jtag_master_master_waitrequest                     => jtag_master_master_waitrequest,                                --                                             .waitrequest
			jtag_master_master_byteenable                      => jtag_master_master_byteenable,                                 --                                             .byteenable
			jtag_master_master_read                            => jtag_master_master_read,                                       --                                             .read
			jtag_master_master_readdata                        => jtag_master_master_readdata,                                   --                                             .readdata
			jtag_master_master_readdatavalid                   => jtag_master_master_readdatavalid,                              --                                             .readdatavalid
			jtag_master_master_write                           => jtag_master_master_write,                                      --                                             .write
			jtag_master_master_writedata                       => jtag_master_master_writedata,                                  --                                             .writedata
			mm_bridge_m0_address                               => mm_bridge_m0_address,                                          --                                 mm_bridge_m0.address
			mm_bridge_m0_waitrequest                           => mm_bridge_m0_waitrequest,                                      --                                             .waitrequest
			mm_bridge_m0_burstcount                            => mm_bridge_m0_burstcount,                                       --                                             .burstcount
			mm_bridge_m0_byteenable                            => mm_bridge_m0_byteenable,                                       --                                             .byteenable
			mm_bridge_m0_read                                  => mm_bridge_m0_read,                                             --                                             .read
			mm_bridge_m0_readdata                              => mm_bridge_m0_readdata,                                         --                                             .readdata
			mm_bridge_m0_readdatavalid                         => mm_bridge_m0_readdatavalid,                                    --                                             .readdatavalid
			mm_bridge_m0_write                                 => mm_bridge_m0_write,                                            --                                             .write
			mm_bridge_m0_writedata                             => mm_bridge_m0_writedata,                                        --                                             .writedata
			mm_bridge_m0_debugaccess                           => mm_bridge_m0_debugaccess,                                      --                                             .debugaccess
			vga_dma_avalon_dma_master_address                  => vga_dma_avalon_dma_master_address,                             --                    vga_dma_avalon_dma_master.address
			vga_dma_avalon_dma_master_waitrequest              => vga_dma_avalon_dma_master_waitrequest,                         --                                             .waitrequest
			vga_dma_avalon_dma_master_read                     => vga_dma_avalon_dma_master_read,                                --                                             .read
			vga_dma_avalon_dma_master_readdata                 => vga_dma_avalon_dma_master_readdata,                            --                                             .readdata
			vga_dma_avalon_dma_master_readdatavalid            => vga_dma_avalon_dma_master_readdatavalid,                       --                                             .readdatavalid
			vga_dma_avalon_dma_master_lock                     => vga_dma_avalon_dma_master_lock,                                --                                             .lock
			key_s1_address                                     => mm_interconnect_0_key_s1_address,                              --                                       key_s1.address
			key_s1_write                                       => mm_interconnect_0_key_s1_write,                                --                                             .write
			key_s1_readdata                                    => mm_interconnect_0_key_s1_readdata,                             --                                             .readdata
			key_s1_writedata                                   => mm_interconnect_0_key_s1_writedata,                            --                                             .writedata
			key_s1_chipselect                                  => mm_interconnect_0_key_s1_chipselect,                           --                                             .chipselect
			led_r_s1_address                                   => mm_interconnect_0_led_r_s1_address,                            --                                     led_r_s1.address
			led_r_s1_write                                     => mm_interconnect_0_led_r_s1_write,                              --                                             .write
			led_r_s1_readdata                                  => mm_interconnect_0_led_r_s1_readdata,                           --                                             .readdata
			led_r_s1_writedata                                 => mm_interconnect_0_led_r_s1_writedata,                          --                                             .writedata
			led_r_s1_chipselect                                => mm_interconnect_0_led_r_s1_chipselect,                         --                                             .chipselect
			leg_g_s1_address                                   => mm_interconnect_0_leg_g_s1_address,                            --                                     leg_g_s1.address
			leg_g_s1_write                                     => mm_interconnect_0_leg_g_s1_write,                              --                                             .write
			leg_g_s1_readdata                                  => mm_interconnect_0_leg_g_s1_readdata,                           --                                             .readdata
			leg_g_s1_writedata                                 => mm_interconnect_0_leg_g_s1_writedata,                          --                                             .writedata
			leg_g_s1_chipselect                                => mm_interconnect_0_leg_g_s1_chipselect,                         --                                             .chipselect
			ps2_avalon_ps2_slave_address                       => mm_interconnect_0_ps2_avalon_ps2_slave_address,                --                         ps2_avalon_ps2_slave.address
			ps2_avalon_ps2_slave_write                         => mm_interconnect_0_ps2_avalon_ps2_slave_write,                  --                                             .write
			ps2_avalon_ps2_slave_read                          => mm_interconnect_0_ps2_avalon_ps2_slave_read,                   --                                             .read
			ps2_avalon_ps2_slave_readdata                      => mm_interconnect_0_ps2_avalon_ps2_slave_readdata,               --                                             .readdata
			ps2_avalon_ps2_slave_writedata                     => mm_interconnect_0_ps2_avalon_ps2_slave_writedata,              --                                             .writedata
			ps2_avalon_ps2_slave_byteenable                    => mm_interconnect_0_ps2_avalon_ps2_slave_byteenable,             --                                             .byteenable
			ps2_avalon_ps2_slave_waitrequest                   => mm_interconnect_0_ps2_avalon_ps2_slave_waitrequest,            --                                             .waitrequest
			ps2_avalon_ps2_slave_chipselect                    => mm_interconnect_0_ps2_avalon_ps2_slave_chipselect,             --                                             .chipselect
			sdram_controller_s1_address                        => mm_interconnect_0_sdram_controller_s1_address,                 --                          sdram_controller_s1.address
			sdram_controller_s1_write                          => mm_interconnect_0_sdram_controller_s1_write,                   --                                             .write
			sdram_controller_s1_read                           => mm_interconnect_0_sdram_controller_s1_read,                    --                                             .read
			sdram_controller_s1_readdata                       => mm_interconnect_0_sdram_controller_s1_readdata,                --                                             .readdata
			sdram_controller_s1_writedata                      => mm_interconnect_0_sdram_controller_s1_writedata,               --                                             .writedata
			sdram_controller_s1_byteenable                     => mm_interconnect_0_sdram_controller_s1_byteenable,              --                                             .byteenable
			sdram_controller_s1_readdatavalid                  => mm_interconnect_0_sdram_controller_s1_readdatavalid,           --                                             .readdatavalid
			sdram_controller_s1_waitrequest                    => mm_interconnect_0_sdram_controller_s1_waitrequest,             --                                             .waitrequest
			sdram_controller_s1_chipselect                     => mm_interconnect_0_sdram_controller_s1_chipselect,              --                                             .chipselect
			sev_seg03_s1_address                               => mm_interconnect_0_sev_seg03_s1_address,                        --                                 sev_seg03_s1.address
			sev_seg03_s1_write                                 => mm_interconnect_0_sev_seg03_s1_write,                          --                                             .write
			sev_seg03_s1_readdata                              => mm_interconnect_0_sev_seg03_s1_readdata,                       --                                             .readdata
			sev_seg03_s1_writedata                             => mm_interconnect_0_sev_seg03_s1_writedata,                      --                                             .writedata
			sev_seg03_s1_chipselect                            => mm_interconnect_0_sev_seg03_s1_chipselect,                     --                                             .chipselect
			sev_seg47_s1_address                               => mm_interconnect_0_sev_seg47_s1_address,                        --                                 sev_seg47_s1.address
			sev_seg47_s1_write                                 => mm_interconnect_0_sev_seg47_s1_write,                          --                                             .write
			sev_seg47_s1_readdata                              => mm_interconnect_0_sev_seg47_s1_readdata,                       --                                             .readdata
			sev_seg47_s1_writedata                             => mm_interconnect_0_sev_seg47_s1_writedata,                      --                                             .writedata
			sev_seg47_s1_chipselect                            => mm_interconnect_0_sev_seg47_s1_chipselect,                     --                                             .chipselect
			sram_0_avalon_sram_slave_address                   => mm_interconnect_0_sram_0_avalon_sram_slave_address,            --                     sram_0_avalon_sram_slave.address
			sram_0_avalon_sram_slave_write                     => mm_interconnect_0_sram_0_avalon_sram_slave_write,              --                                             .write
			sram_0_avalon_sram_slave_read                      => mm_interconnect_0_sram_0_avalon_sram_slave_read,               --                                             .read
			sram_0_avalon_sram_slave_readdata                  => mm_interconnect_0_sram_0_avalon_sram_slave_readdata,           --                                             .readdata
			sram_0_avalon_sram_slave_writedata                 => mm_interconnect_0_sram_0_avalon_sram_slave_writedata,          --                                             .writedata
			sram_0_avalon_sram_slave_byteenable                => mm_interconnect_0_sram_0_avalon_sram_slave_byteenable,         --                                             .byteenable
			sram_0_avalon_sram_slave_readdatavalid             => mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid,      --                                             .readdatavalid
			switch_s1_address                                  => mm_interconnect_0_switch_s1_address,                           --                                    switch_s1.address
			switch_s1_write                                    => mm_interconnect_0_switch_s1_write,                             --                                             .write
			switch_s1_readdata                                 => mm_interconnect_0_switch_s1_readdata,                          --                                             .readdata
			switch_s1_writedata                                => mm_interconnect_0_switch_s1_writedata,                         --                                             .writedata
			switch_s1_chipselect                               => mm_interconnect_0_switch_s1_chipselect,                        --                                             .chipselect
			vga_dma_avalon_dma_control_slave_address           => mm_interconnect_0_vga_dma_avalon_dma_control_slave_address,    --             vga_dma_avalon_dma_control_slave.address
			vga_dma_avalon_dma_control_slave_write             => mm_interconnect_0_vga_dma_avalon_dma_control_slave_write,      --                                             .write
			vga_dma_avalon_dma_control_slave_read              => mm_interconnect_0_vga_dma_avalon_dma_control_slave_read,       --                                             .read
			vga_dma_avalon_dma_control_slave_readdata          => mm_interconnect_0_vga_dma_avalon_dma_control_slave_readdata,   --                                             .readdata
			vga_dma_avalon_dma_control_slave_writedata         => mm_interconnect_0_vga_dma_avalon_dma_control_slave_writedata,  --                                             .writedata
			vga_dma_avalon_dma_control_slave_byteenable        => mm_interconnect_0_vga_dma_avalon_dma_control_slave_byteenable  --                                             .byteenable
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => sdram_pll_reset_source_reset,   -- reset_in0.reset
			clk            => sdram_pll_sys_clk_clk,          --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => jtag_master_master_reset_reset,     -- reset_in0.reset
			clk            => sdram_pll_sys_clk_clk,              --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_003 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => vga_pll_reset_source_reset,         -- reset_in0.reset
			clk            => vga_pll_vga_clk_clk,                --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_sdram_controller_s1_read_ports_inv <= not mm_interconnect_0_sdram_controller_s1_read;

	mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_controller_s1_byteenable;

	mm_interconnect_0_sdram_controller_s1_write_ports_inv <= not mm_interconnect_0_sdram_controller_s1_write;

	mm_interconnect_0_leg_g_s1_write_ports_inv <= not mm_interconnect_0_leg_g_s1_write;

	mm_interconnect_0_switch_s1_write_ports_inv <= not mm_interconnect_0_switch_s1_write;

	mm_interconnect_0_key_s1_write_ports_inv <= not mm_interconnect_0_key_s1_write;

	mm_interconnect_0_led_r_s1_write_ports_inv <= not mm_interconnect_0_led_r_s1_write;

	mm_interconnect_0_sev_seg03_s1_write_ports_inv <= not mm_interconnect_0_sev_seg03_s1_write;

	mm_interconnect_0_sev_seg47_s1_write_ports_inv <= not mm_interconnect_0_sev_seg47_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of AvalonMM
